* C:\Users\hp\eSim-Workspace\CM\CM.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 11/08/24 23:22:27

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_I1-Pad2_ GND Net-_X1-Pad3_ Net-_SC1-Pad1_ Net-_SC1-Pad2_ GND avsd_opamp		
X2  Net-_U2-Pad1_ GND Net-_SC2-Pad1_ Net-_X1-Pad3_ Net-_SC3-Pad2_ GND avsd_opamp		
I1  Net-_I1-Pad1_ Net-_I1-Pad2_ dc		
U1  Net-_SC4-Pad1_ Net-_SC1-Pad1_ plot_i2		
v3  Net-_U2-Pad1_ GND DC		
v1  Net-_X1-Pad3_ GND DC		
v2  Net-_I1-Pad2_ GND DC		
U2  Net-_U2-Pad1_ Net-_SC3-Pad1_ plot_i2		
scmode1  SKY130mode		
SC3  Net-_SC3-Pad1_ Net-_SC3-Pad2_ Net-_SC2-Pad1_ Net-_SC2-Pad1_ sky130_fd_pr__nfet_01v8		
SC2  Net-_SC2-Pad1_ Net-_SC1-Pad2_ GND GND sky130_fd_pr__nfet_01v8		
SC1  Net-_SC1-Pad1_ Net-_SC1-Pad2_ GND GND sky130_fd_pr__nfet_01v8		
SC4  Net-_SC4-Pad1_ Net-_I1-Pad1_ ? sky130_fd_pr__res_high_po_0p69		

.end
