* C:\Users\hp\eSim-Workspace\CM\CM.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 11/08/24 20:12:33

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X1  Net-_I1-Pad2_ GND Net-_X1-Pad3_ Net-_M1-Pad1_ Net-_M1-Pad2_ GND avsd_opamp		
X2  Net-_U2-Pad1_ GND Net-_M2-Pad1_ Net-_X1-Pad3_ Net-_M3-Pad2_ GND avsd_opamp		
I1  Net-_I1-Pad1_ Net-_I1-Pad2_ dc		
U1  Net-_I1-Pad1_ Net-_M1-Pad1_ plot_i2		
v3  Net-_U2-Pad1_ GND DC		
v1  Net-_X1-Pad3_ GND DC		
v2  Net-_I1-Pad2_ GND DC		
U2  Net-_U2-Pad1_ Net-_M3-Pad1_ plot_i2		
M3  Net-_M3-Pad1_ Net-_M3-Pad2_ Net-_M2-Pad1_ Net-_M2-Pad1_ eSim_MOS_N		
M1  Net-_M1-Pad1_ Net-_M1-Pad2_ GND GND eSim_MOS_N		
M2  Net-_M2-Pad1_ Net-_M1-Pad2_ GND GND eSim_MOS_N		
scmode1  SKY130mode		

.end
